module gaussian_blur;
    // Parameters for image dimensions and kernel size
    parameter integer IMG_WIDTH = 247;  // Width of the image (modify as needed)
    parameter integer IMG_HEIGHT = 242; // Height of the image (modify as needed)
    parameter integer KERNEL_SIZE = 9;  // Gaussian kernel size (NxN, modify as needed)

    // Gaussian kernel coefficients - dynamically generated based on KERNEL_SIZE
    real GAUSSIAN_KERNEL[0:KERNEL_SIZE-1][0:KERNEL_SIZE-1];

    // File handles
    integer input_file, output_file;
    integer i, j, m, n, idx;

    // Memory to hold the image and result
    reg [7:0] image[0:IMG_HEIGHT-1][0:IMG_WIDTH-1];
    real blurred_image[0:IMG_HEIGHT-1][0:IMG_WIDTH-1];

    // Temporary storage for pixel value and sum
    real pixel_sum;
    reg [7:0] temp_pixel;

    // Variables for Gaussian kernel generation
    real sigma;
    real sum;

    initial begin
        // Initialize Gaussian kernel variables
        sigma = KERNEL_SIZE / 6.0; // Standard deviation approximation
        sum = 0.0;

        // Generate Gaussian kernel dynamically based on KERNEL_SIZE
        for (m = 0; m < KERNEL_SIZE; m = m + 1) begin
            for (n = 0; n < KERNEL_SIZE; n = n + 1) begin
                GAUSSIAN_KERNEL[m][n] = $exp(-((m-KERNEL_SIZE/2)*(m-KERNEL_SIZE/2) + (n-KERNEL_SIZE/2)*(n-KERNEL_SIZE/2)) / (2*sigma*sigma));
                sum = sum + GAUSSIAN_KERNEL[m][n];
            end
        end
        // Normalize the kernel
        for (m = 0; m < KERNEL_SIZE; m = m + 1) begin
            for (n = 0; n < KERNEL_SIZE; n = n + 1) begin
                GAUSSIAN_KERNEL[m][n] = GAUSSIAN_KERNEL[m][n] / sum;
            end
        end

        // Open input and output files
        input_file = $fopen("input_image.txt", "r");
        output_file = $fopen("output_image.txt", "w");

        // Check if files are opened successfully
        if (input_file == 0) begin
            $display("Error: Cannot open input_image.txt");
            $finish;
        end

        if (output_file == 0) begin
            $display("Error: Cannot open output_image.txt");
            $finish;
        end

        // Read the input image into memory
        for (i = 0; i < IMG_HEIGHT; i = i + 1) begin
            for (j = 0; j < IMG_WIDTH; j = j + 1) begin
                idx = $fscanf(input_file, "%d", temp_pixel);
                image[i][j] = temp_pixel;
            end
        end

        // Apply Gaussian blur
        for (i = KERNEL_SIZE/2; i < IMG_HEIGHT-KERNEL_SIZE/2; i = i + 1) begin
            for (j = KERNEL_SIZE/2; j < IMG_WIDTH-KERNEL_SIZE/2; j = j + 1) begin
                pixel_sum = 0.0;
                // Convolve with the Gaussian kernel
                for (m = 0; m < KERNEL_SIZE; m = m + 1) begin
                    for (n = 0; n < KERNEL_SIZE; n = n + 1) begin
                        pixel_sum = pixel_sum + image[i+m-KERNEL_SIZE/2][j+n-KERNEL_SIZE/2] * GAUSSIAN_KERNEL[m][n];
                    end
                end
                // Store the blurred value
                blurred_image[i][j] = pixel_sum;
            end
        end

        // Write the blurred image to the output file
        for (i = 0; i < IMG_HEIGHT; i = i + 1) begin
            for (j = 0; j < IMG_WIDTH; j = j + 1) begin
                $fwrite(output_file, "%d", $rtoi(blurred_image[i][j]));
                if (j < IMG_WIDTH-1) $fwrite(output_file, " "); // Add space between pixels
            end
            $fwrite(output_file, "\n"); // Add a newline at the end of each row
        end

        // Close the files
        $fclose(input_file);
        $fclose(output_file);

        $display("Gaussian blur completed. Output written to output_image.txt");
        $finish;
    end
endmodule
